module DataMemoryUnit(
    input wire clk,
    input wire memWrite,
    input wire memRead,
    input wire [31:0] address,
    input wire [31:0] writeData,
    output reg [31:0] readData,
    output wire [31:0] memory8, memory12, memory16, memory20
);

    reg [31:0] memory [0:1023];

    initial begin
        memory[0] = 8'b00000000;
        memory[1] = 8'b00000000;
        memory[2] = 8'b00000000;
        memory[3] = 8'b00000000;     // dummy
        //000000 00000 00000 00000 00000 000000   
        memory[4] = 8'b00100001;
        memory[5] = 8'b00001000;
        memory[6] = 8'b00000000;
        memory[7] = 8'b00001000;     // addi $t0, $t0, 8
        //001000 01000 01000 0000000000001000
        memory[8] = 8'b00100001;
        memory[9] = 8'b00101001;
        memory[10] = 8'b00000000;
        memory[11] = 8'b00001000;     // addi $t1, $t1, 8
        //001000 01001 01001 0000000000001000    
        memory[12] = 8'b00010001;
        memory[13] = 8'b00001001;
        memory[14] = 8'b00000000;
        memory[15] = 8'b01100100;     // beq $t0, $t1, 100
        //000100 01000 01001 0000000001100100
        memory[16] = 8'b00000001;
        memory[17] = 8'b00101000;
        memory[18] = 8'b01011000;
        memory[19] = 8'b00100000;    // add $t3, $t1, $t0
        //000000 01001 01000 01011 00000 100000
        memory[20] = 8'b00000001;
        memory[21] = 8'b00101001;
        memory[22] = 8'b01011000;
        memory[23] = 8'b00100000;    // add $t3, $t1, $t1
        //000000 01001 01001 01011 00000 100000
        memory[416] = 8'b00000001;
        memory[417] = 8'b00101000;
        memory[418] = 8'b01010000;
        memory[419] = 8'b00100000;   // add $t2, $t1, $t0
        //000000 01001 01000 01010 00000 100000
        memory[420] = 8'b00100001;
        memory[421] = 8'b00001000;
        memory[422] = 8'b00000000;
        memory[423] = 8'b00001111;       // addi $t0, $t0, 15
        //001000 01000 01000 0000000000001000
        memory[424] = 8'b00100001;
        memory[425] = 8'b00101001;
        memory[426] = 8'b00000000;
        memory[427] = 8'b00000101;       // addi $t1, $t1, 5
        //001000 01001 01001 0000000000001000  
        memory[428] = 8'b00000001;
        memory[429] = 8'b00101000;
        memory[430] = 8'b01010000;
        memory[431] = 8'b00101010;      // slt $t2, $t1, $t0
        //000000 01001 01000 01010 00000 101010
        
/*
        memory[0] = 8'b00000000;
        memory[1] = 8'b00000000;
        memory[2] = 8'b00000000;
        memory[3] = 8'b00000000;     // dummy
        //000000 00000 00000 00000 00000 000000        
        memory[4] = 8'b00100001;
        memory[5] = 8'b00001000;
        memory[6] = 8'b00000000;
        memory[7] = 8'b00000000;     // addi $t0, $t0, 0
        //001000 01000 01000 0000000000000000
        memory[8] = 8'b00100001;
        memory[9] = 8'b00101001;
        memory[10] = 8'b00000000;
        memory[11] = 8'b00000001;     // addi $t1, $t1, 1
        //001000 01001 01001 0000000000000001        
        memory[12] = 8'b00000001;
        memory[13] = 8'b00001001;
        memory[14] = 8'b01010000;
        memory[15] = 8'b00100100;    // and $t2, $t0, $t1
        //000000 01000 01001 01010 00000 100100
        memory[16] = 8'b00000001;
        memory[17] = 8'b00001001;
        memory[18] = 8'b01011000;
        memory[19] = 8'b00100101;    // or $t3, $t0, $t1
        //000000 01000 01001 01011 00000 100101
        memory[20] = 8'b00000001;
        memory[21] = 8'b00101001;
        memory[22] = 8'b01010000;
        memory[23] = 8'b00100100;    // and $t2, $t1, $t1
        //000000 01001 01001 01010 00000 100100
        memory[24] = 8'b00000001;
        memory[25] = 8'b00001000;
        memory[26] = 8'b01011000;
        memory[27] = 8'b00100101;    // or $t3, $t0, $t0
        //000000 01000 01000 01011 00000 100101
        memory[28] = 8'b00000001;
        memory[29] = 8'b00001001;
        memory[30] = 8'b01000000;
        memory[31] = 8'b00101010;    // slt $t0, $t0, $t1
        //000000 01000 01001 01000 00000 101010
        memory[32] = 8'b00000001;
        memory[33] = 8'b00001001;
        memory[34] = 8'b01011000;
        memory[35] = 8'b00100100;    // and $t3, $t0, $t1
        //000000 01000 01001 01011 00000 100100
        memory[36] = 8'b00000001;
        memory[37] = 8'b00101000;
        memory[38] = 8'b01010000;
        memory[39] = 8'b00100000;    // add $t2, $t1, $t0
        //000000 01001 01000 01010 00000 100000
        memory[40] = 8'b00000001;
        memory[41] = 8'b01001001;
        memory[42] = 8'b01011000;
        memory[43] = 8'b00100000;    // add $t3, $t2, $t1
        //000000 01010 01001 01011 00000 100000
        memory[44] = 8'b00000001;
        memory[45] = 8'b01101001;
        memory[46] = 8'b01011000;
        memory[47] = 8'b00100010;    // sub $t3, $t3, $t1
        //000000 01011 01001 01011 00000 100010
        memory[48] = 8'b10001101;
        memory[49] = 8'b00001001;
        memory[50] = 8'b00000000;
        memory[51] = 8'b00000111;    // lw $t1, 7($t0)
        //100011 01000 01001 00000000000111
        memory[52] = 8'b00000001;
        memory[53] = 8'b00101010;
        memory[54] = 8'b01000000;
        memory[55] = 8'b00100010;    // sub $t0, $t1, $t2
        //000000 01001 01010 01000 00000 100010
        memory[56] = 8'b10101101;
        memory[57] = 8'b00001000;
        memory[58] = 8'b00000000;
        memory[59] = 8'b00000110;    // sw $t0, 6($t0)
        //101011 01000 01000 0000000000000101 
*/
    always @(negedge clk) begin
        if (memWrite)
            memory[address] <= writeData;
        if (memRead)
            readData <= memory[address];
    end
    
    assign memory8 = memory[8];
    assign memory12 = memory[12];
    assign memory16 = memory[16];
    assign memory20 = memory[20];

endmodule
